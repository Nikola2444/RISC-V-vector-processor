
 `define DDR_DEPTH 4096

