//`define CONV_1X1

`define PD_SIZE 1
`define FR_SIZE 3
`define IM_SIZE 56
`define IN_D    64
`define OUT_D   64
`define INSTR_MEM_SIZE
`define DDR_DEPTH 1500000
`define V_LANES  8
`define VLEN  4096
`define VRF_DEPTH `VLEN/`V_LANES
