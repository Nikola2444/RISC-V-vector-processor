`define CONV_1X1

`define PD_SIZE 1
`define FR_SIZE 1
`define IM_SIZE 3
`define IN_D    512
`define OUT_D   16
`define INSTR_MEM_SIZE
`define DDR_DEPTH 1500000
`define V_LANES  8
`define VLEN  4096
`define VRF_DEPTH `VLEN/`V_LANES
