
`define DDR_DEPTH 8192*4
`define V_LANES  4
`define VLEN  4096
`define VRF_DEPTH `VLEN/`V_LANES
